// HDLBits: Hello, World (wire)
module hello_wire(input a, output b);
  assign b = a;
endmodule
